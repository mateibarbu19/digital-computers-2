module test_ram();

endmodule
 
