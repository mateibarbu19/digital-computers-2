../lab-08/defines.vh